/* Autor: Sergio Garino Vargas
 * Carné: B73157
 * Fecha de entrega: 9/12/2022
 */


 module PARITY_SEVEN ( input [6:0] x_n,
                       output R);

    

 endmodule